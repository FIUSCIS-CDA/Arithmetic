///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: SESL
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020, 2025 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbenchSESL();
`include "../Test/Test.v"


//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing SESL16_32
reg[15:0] A_16;
wire[31:0] A_32;
SESL16_32 mySESL16(.A(A_16), .Y(A_32));
//////////////////////////////////////////////////////////////////////////////////////////////////////


initial begin 
////////////////////////////////////////////////////////////////////////////////////////
// Test: 114 (16 to 32)
$display("Testing: 114");
A_16=114; #10;
verifyEqual32(A_32, 114*4);
////////////////////////////////////////////////////////////////////////////////////////
 
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule
