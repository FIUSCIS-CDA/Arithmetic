///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: INC4_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020, 2025 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbenchINC4();
`include "../Test/Test.v"


//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing INC4
// Also tests Adder_32
reg[31:0] A;
wire[31:0] Result;
wire overflow;
INC4_32 myINC4(.A(A), .Overflow(overflow), .S(Result));
//////////////////////////////////////////////////////////////////////////////////////////////////////

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 + 4 = 49
$display("Testing: 45 + 4 = 49");
A=45;    #10; 
verifyEqual32(Result, 49);
$display("  Ensuring no overflow"); 
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule
