///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: ALU_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020, 2025 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbenchALU();
`include "../Test/Test.v"


//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing the ALU will test:
// ALU_32
// AND_32
// Adder_32
// Less_32
// Log2_32
// Multiplier_32
// NOT_32 (in Subtractor_32)
// OR_32
// OneBitAdder (in Adder_32)
// OneBitAdderHalf (in Multiplier_32)
// SLL_32
// ZE5_32 (in ALU_32)
reg[31:0] A;
reg[31:0] B;
reg[4:0] H;
reg[2:0] alu_op; 
wire[31:0] Result;
wire overflow;
ALU_32 myALU(.A(A), .alu_op(alu_op), .B(B), .H(H),  .Overflow(overflow), .Result(Result));
//////////////////////////////////////////////////////////////////////////////////////////////////////

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 & 21 = 5
$display("Testing: 45 & 21 = 5");
A=45; alu_op=3'b000; B=21;   #10; 
verifyEqual32(Result, A&B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 | 21 = 61
$display("Testing: 45 | 21 = 61");
A=45; alu_op=3'b001; B=21;   #10; 
verifyEqual32(Result, A|B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 + 21 = 66
$display("Testing: 45 + 21 = 66");
A=45; alu_op=3'b010; B=21;   #10; 
verifyEqual32(Result, A+B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0); 
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 - 21 = 24
$display("Testing: 45 - 21 = 24");
A=45; alu_op=3'b011; B=21;   #10; 
verifyEqual32(Result, A-B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 < 21 = 0
$display("Testing: 45 < 21 = 0");
A=45; alu_op=3'b100; B=21;   #10; 
verifyEqual32(Result, A<B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 21 < 45 = 1
$display("Testing: 21 < 45 = 0");
A=21; alu_op=3'b100; B=45;   #10; 
verifyEqual32(Result, A<B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////


////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)+1 overflows
$display("Testing if (2^31-1)+1 overflows: 1");
A = 2147483647; B = 1; alu_op=3'b010; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)+(-1) overflows
$display("Testing if (-2^31)+(-1) overflows: 1");
A = -2147483648; B = -1; alu_op=3'b010; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)-1 overflows
$display("Testing if (-2^31)-1 overflows: 1");
A = -2147483648; B = 1; alu_op=3'b011; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)-(-1) overflows
$display("Testing if (2^31-1)-(-1) overflows: 1");
A = 2147483647; B = -1; alu_op=3'b011; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)<(-1) overflows (it will, < uses -)
$display("Testing if (2^31-1)<(-1) overflows: 1");
A = 2147483647; B = -1; alu_op=3'b100; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)<(1) overflows (it will, < uses -)
$display("Testing if (-2^31)<(1) overflows: 1");
A = -2147483648; B = 1; alu_op=3'b100; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 * 2 = 90
$display("Testing: 45 * 2 = 90");
A=45; B=2; alu_op=3'b101;   #10; 
verifyEqual32(Result, A*B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 << 2 = 180
$display("Testing: 45 << 2 = 180");
B=45; H=2; alu_op=3'b110;   #10; 
verifyEqual32(Result, B*4);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(32) = 5
$display("Testing: log2(32) = 5");
A=32; alu_op=3'b111;   #10; 
verifyEqual32(Result, 5);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule
