///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: EQ
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020, 2025 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbenchEQ();
`include "../Test/Test.v"


//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing EQ_32
reg[31:0] A_32;
reg[31:0] B_32;
wire isEqual_32;
EQ_32 myEQ32(.A(A_32), .B(B_32), .Y(isEqual_32));
//////////////////////////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////////////////////////
// Testing EQ_NONZERO_5
reg[4:0] A_5;
reg[4:0] B_5;
wire isEqual_5;
EQ_NONZERO_5 myEQNZ5(.reg1(A_5), .reg2(B_5), .Y(isEqual_5));
//////////////////////////////////////////////////////////////////////////////////////////////////////

initial begin 
////////////////////////////////////////////////////////////////////////////////////////
// Test: 5 == 5 (True)
$display("Testing: 5 == 5 (True)");
A_32=5; B_32=5;   #10; 
verifyEqual32(isEqual_32, 1);
// Test: 5 == 7 (False)
$display("Testing: 5 == 7 (False)");
A_32=5; B_32=7;   #10; 
verifyEqual32(isEqual_32, 0);
// Test: 5 == 5 (True)
$display("Testing: 5 == 5 (True)");
A_5=5; B_5=5;   #10; 
verifyEqual32(isEqual_5, 1);
// Test: 5 == 0 (False)
$display("Testing: 5 == 0 (False)");
A_5=5; B_5=0;   #10; 
verifyEqual5(isEqual_5, 0);
// Test: 0 == 0 (False, inputs are zero)
$display("Testing: 0 == 0 (False)");
A_5=0; B_5=0;   #10; 
verifyEqual5(isEqual_5, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule
